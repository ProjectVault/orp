0: wb_sdhc_dat_o <= 32'heb3c906d;
1: wb_sdhc_dat_o <= 32'h6b66732e;
2: wb_sdhc_dat_o <= 32'h66617400;
3: wb_sdhc_dat_o <= 32'h02010100;
4: wb_sdhc_dat_o <= 32'h01000200;
5: wb_sdhc_dat_o <= 32'h08f80600;
6: wb_sdhc_dat_o <= 32'h3f00ff00;
9: wb_sdhc_dat_o <= 32'h800029f9;
10: wb_sdhc_dat_o <= 32'h39c5584e;
11: wb_sdhc_dat_o <= 32'h4f204e41;
12: wb_sdhc_dat_o <= 32'h4d452020;
13: wb_sdhc_dat_o <= 32'h20204641;
14: wb_sdhc_dat_o <= 32'h54313220;
15: wb_sdhc_dat_o <= 32'h20200e1f;
16: wb_sdhc_dat_o <= 32'hbe5b7cac;
17: wb_sdhc_dat_o <= 32'h22c0740b;
18: wb_sdhc_dat_o <= 32'h56b40ebb;
19: wb_sdhc_dat_o <= 32'h0700cd10;
20: wb_sdhc_dat_o <= 32'h5eebf032;
21: wb_sdhc_dat_o <= 32'he4cd16cd;
22: wb_sdhc_dat_o <= 32'h19ebfe54;
23: wb_sdhc_dat_o <= 32'h68697320;
24: wb_sdhc_dat_o <= 32'h6973206e;
25: wb_sdhc_dat_o <= 32'h6f742061;
26: wb_sdhc_dat_o <= 32'h20626f6f;
27: wb_sdhc_dat_o <= 32'h7461626c;
28: wb_sdhc_dat_o <= 32'h65206469;
29: wb_sdhc_dat_o <= 32'h736b2e20;
30: wb_sdhc_dat_o <= 32'h20506c65;
31: wb_sdhc_dat_o <= 32'h61736520;
32: wb_sdhc_dat_o <= 32'h696e7365;
33: wb_sdhc_dat_o <= 32'h72742061;
34: wb_sdhc_dat_o <= 32'h20626f6f;
35: wb_sdhc_dat_o <= 32'h7461626c;
36: wb_sdhc_dat_o <= 32'h6520666c;
37: wb_sdhc_dat_o <= 32'h6f707079;
38: wb_sdhc_dat_o <= 32'h20616e64;
39: wb_sdhc_dat_o <= 32'h0d0a7072;
40: wb_sdhc_dat_o <= 32'h65737320;
41: wb_sdhc_dat_o <= 32'h616e7920;
42: wb_sdhc_dat_o <= 32'h6b657920;
43: wb_sdhc_dat_o <= 32'h746f2074;
44: wb_sdhc_dat_o <= 32'h72792061;
45: wb_sdhc_dat_o <= 32'h6761696e;
46: wb_sdhc_dat_o <= 32'h202e2e2e;
47: wb_sdhc_dat_o <= 32'h200d0a00;
127: wb_sdhc_dat_o <= 32'h000055aa;
128: wb_sdhc_dat_o <= 32'hf8ffff00;
129: wb_sdhc_dat_o <= 32'h40000560;
130: wb_sdhc_dat_o <= 32'h00ff8f00;
131: wb_sdhc_dat_o <= 32'h09a000ff;
132: wb_sdhc_dat_o <= 32'h0f000000;
896: wb_sdhc_dat_o <= 32'h5246494c;
897: wb_sdhc_dat_o <= 32'h45202020;
898: wb_sdhc_dat_o <= 32'h20202020;
899: wb_sdhc_dat_o <= 32'h0000302c;
900: wb_sdhc_dat_o <= 32'h53465346;
901: wb_sdhc_dat_o <= 32'h0000302c;
902: wb_sdhc_dat_o <= 32'h53460300;
903: wb_sdhc_dat_o <= 32'h00080000;
904: wb_sdhc_dat_o <= 32'h5746494c;
905: wb_sdhc_dat_o <= 32'h45202020;
906: wb_sdhc_dat_o <= 32'h20202020;
907: wb_sdhc_dat_o <= 32'h0000332c;
908: wb_sdhc_dat_o <= 32'h53465346;
909: wb_sdhc_dat_o <= 32'h0000332c;
910: wb_sdhc_dat_o <= 32'h53460700;
911: wb_sdhc_dat_o <= 32'h00080000;
