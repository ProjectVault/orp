0: wb_dat_o <= 32'h18609100;
1: wb_dat_o <= 32'h9c8000ff;
2: wb_dat_o <= 32'hd8032000;
3: wb_dat_o <= 32'hd8032001;
4: wb_dat_o <= 32'h18e00010;
5: wb_dat_o <= 32'ha8e70000;
6: wb_dat_o <= 32'h9c800000;
7: wb_dat_o <= 32'hd8032000;
8: wb_dat_o <= 32'h18c00000;
9: wb_dat_o <= 32'h9cc60001;
10: wb_dat_o <= 32'he4063800;
11: wb_dat_o <= 32'h0ffffffe;
12: wb_dat_o <= 32'h15000000;
13: wb_dat_o <= 32'h9c8000ff;
14: wb_dat_o <= 32'hd8032000;
15: wb_dat_o <= 32'h18c00000;
16: wb_dat_o <= 32'h9cc60001;
17: wb_dat_o <= 32'he4063800;
18: wb_dat_o <= 32'h0ffffffe;
19: wb_dat_o <= 32'h15000000;
20: wb_dat_o <= 32'h03fffff2;
21: wb_dat_o <= 32'h15000000;
