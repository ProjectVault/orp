110: wb_sdhc_dat_o <= 32'h1e03b615;
111: wb_sdhc_dat_o <= 32'h00000020;
112: wb_sdhc_dat_o <= 32'h21000641;
113: wb_sdhc_dat_o <= 32'h01000008;
114: wb_sdhc_dat_o <= 32'h00000008;
127: wb_sdhc_dat_o <= 32'h000055aa;
